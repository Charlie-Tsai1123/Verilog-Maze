module Maze(
    input Clk,
    input Reset,
    input right,
    input left,
    input forward,
    input backward,
    output [7:0] dotrow,
    output [15:0] dotcol,
    output [6:0]out_decimal,
    output [6:0]out,
    output [6:0]win_decimal,
    output [6:0]win
);

wire [127:0] maze_origin;
wire [127:0] maze_with_player;
wire [6:0] player_index;
wire endGame;
wire refresh_maze;

GenerateMaze gen_maze(Clk, refresh_maze, maze_origin);
GetPlayerIndex get_playIdx(Clk, Reset, right, left, forward, backward, maze_origin, refresh_maze, player_index, endGame);
AddPlayer add_player(Clk, player_index, maze_origin, maze_with_player);
DisplayMaze disp_maze(Clk, maze_with_player, dotrow, dotcol);
CountAndGrade count_and_grade(Clk, Reset, endGame, out_decimal, out, win_decimal, win, refresh_maze);
 
endmodule
 
 
module GetPlayerIndex (
    input Clk,
    input Reset,
    input right,
    input left,
    input forward,
    input backward,
    input [127:0] maze,
    input refresh_maze,
    output reg [6:0] id,
    output reg endGame
);
 
reg [31:0] counter = 32'b0;
reg isPressRight = 0;
reg isPressLeft = 0;
reg isPressForward = 0;
reg isPressBackward = 0;
 
initial begin
    id = 7'd126;
end
 
always @(posedge Clk or negedge Reset) begin
    //print the player (maze)
    
    if (!Reset)
    begin
        id <= 7'd126;
        counter <= 32'd0;
        isPressRight <= 0;
        isPressLeft <= 0;
        isPressForward <= 0;
        isPressBackward <= 0;
    end
    else
    begin
        if(counter == 32'd5000) begin
            counter <= 32'b0;
            if(!right && isPressRight == 0) begin
                isPressRight = 1;
                if(maze[id - 7'd1] == 7'd0) begin
                    id <= id - 7'd1;
                end
            end
        
            if(!left && isPressLeft == 0) begin
                isPressLeft = 1;
                if(maze[id + 7'd1] == 7'd0) begin
                    id <= id + 7'd1;
                end
            end
        
            if(!forward && isPressForward == 0) begin
                isPressForward = 1;
                if(maze[id + 7'd16] == 7'd0) begin
                    id <= id + 7'd16;
                end
            end
        
            if(!backward && isPressBackward == 0) begin
                isPressBackward = 1;
                if(maze[id - 7'd16] == 7'd0) begin
                        if(id - 7'd16 == 7'd2) begin
                            id <= 7'd126;
                            endGame <= 1;
                        end else begin
                            id <= id - 7'd16;
                        end
                end
            end
        
            if(right) isPressRight = 0;
            if(left) isPressLeft = 0;
            if(forward) isPressForward = 0;
            if(backward) isPressBackward = 0;
            if(refresh_maze) begin
                id <= 7'd126;
                endGame <= 0;
            end
        end else begin
            counter <= counter + 32'd1; 
        end
    end
    
end
    
endmodule
 
 
module AddPlayer (
    input Clk,
    input [6:0] index,
    input [127:0] maze_in,
    output reg [127:0] maze_out
);
 
reg [31:0] counter;
reg flash;
 
always @(posedge Clk)
begin
    if (counter == 32'd12500000)
    begin
        counter <= 32'd0;
        flash <= ~flash;
        if (flash == 1'b1)
            maze_out <= (maze_in | (128'd1 << index));
        else
            maze_out <= maze_in;
    end
    else
    begin
        counter <= counter + 32'd1;
    end
end
    
endmodule
 
 
module DisplayMaze (
    input Clk,
    input [127:0] maze,
    output reg [7:0] dotrow,
    output reg [15:0] dotcol
);
 
reg [31:0] counter;
reg [2:0] setLight;
 
always @(posedge Clk) begin
        
    //print the player (maze)
    if(counter == 32'd5000)
    begin
        counter <= 32'b0;
        
        if(setLight==3'd7) setLight <= 3'd0;
        else setLight <= setLight+1;
        
        case(setLight)
            3'd7:dotrow<=8'b01111111;
            3'd6:dotrow<=8'b10111111;
            3'd5:dotrow<=8'b11011111;
            3'd4:dotrow<=8'b11101111;
            3'd3:dotrow<=8'b11110111;
            3'd2:dotrow<=8'b11111011;
            3'd1:dotrow<=8'b11111101;
            3'd0:dotrow<=8'b11111110;
        endcase
        
        dotcol[0] <= maze[setLight*16];
        dotcol[1] <= maze[setLight*16 + 1];
        dotcol[2] <= maze[setLight*16 + 2];
        dotcol[3] <= maze[setLight*16 + 3];
        dotcol[4] <= maze[setLight*16 + 4];
        dotcol[5] <= maze[setLight*16 + 5];
        dotcol[6] <= maze[setLight*16 + 6];
        dotcol[7] <= maze[setLight*16 + 7];
        dotcol[8] <= maze[setLight*16 + 8];
        dotcol[9] <= maze[setLight*16 + 9];
        dotcol[10] <= maze[setLight*16 + 10];
        dotcol[11] <= maze[setLight*16 + 11];
        dotcol[12] <= maze[setLight*16 + 12];
        dotcol[13] <= maze[setLight*16 + 13];
        dotcol[14] <= maze[setLight*16 + 14];
        dotcol[15] <= maze[setLight*16 + 15];
    end 
    else counter <= counter + 32'd1; 
end
endmodule
 
 
module GenerateMaze (
    input Clk,
    input refresh_maze,
    output reg [127:0] maze
);
 
reg [31:0] random;
reg [31:0] index;
 
initial begin
    maze = 128'b10111111111111111000000000000011111111111111101110000010000000111011101011111111100010000000001111111111111110111111111111111011;
    random = 32'd0;
end

// random
always @(posedge Clk) 
begin
    if (random == 32'd99)
        random <= 32'd0;
    else
        random <= random + 32'd1;
end

always @(posedge refresh_maze)
begin
    if (refresh_maze) begin
        index <= random;
        case (index)
            32'd0: maze <= 128'b10111111111111111000000000000011111111111111101110000010000000111011101011111111100010000000001111111111111110111111111111111011;
            32'd1: maze <= 128'b10111111111111111000001000100011111110101010101110100010101010111010111010111011100000001000001111111111111110111111111111111011;
            32'd2: maze <= 128'b10111111111111111010000000100011101011111010111110101000101000111010101110111011100010000000001111111111111110111111111111111011;
            32'd3: maze <= 128'b10111111111111111000000000100011111111111011101110000000100010111011101111101011100010000000001111111111111110111111111111111011;
            32'd4: maze <= 128'b10111111111111111000001000100011111110101010101110001010100010111011101111111011100000000000001111111111111110111111111111111011;
            32'd5: maze <= 128'b10111111111111111000000000000011111111111111101110001000100000111011101010111111100000100000001111111111111110111111111111111011;
            32'd6: maze <= 128'b10111111111111111010001000000011101010101111101110101010001000111010101110101111100010000010001111111111111110111111111111111011;
            32'd7: maze <= 128'b10111111111111111010000000000011101011111111101110001000100000111111101010111111100000100000001111111111111110111111111111111011;
            32'd8: maze <= 128'b10111111111111111010001000100011101010101010101110101010101010111010101010111011100010001000001111111111111110111111111111111011;
            32'd9: maze <= 128'b10111111111111111000000010000011111111101011101110001000100010111010101111111011101000000000001111111111111110111111111111111011;
            32'd10: maze <= 128'b10111111111111111010000010000011101011101011101110101010100010111010101011111011100010000000001111111111111110111111111111111011;
            32'd11: maze <= 128'b10111111111111111000001000001011111110101110101110000010100010111011111010111011100000001000001111111111111110111111111111111011;
            32'd12: maze <= 128'b10111111111111111000001000000011111110111011101110000010001010111011111011101011100000001000001111111111111110111111111111111011;
            32'd13: maze <= 128'b10111111111111111000100000000011111010111111101110001010000010111011101010111011100000101000001111111111111110111111111111111011;
            32'd14: maze <= 128'b10111111111111111010000010000011101010101010111110101010101000111011101011111011100000100000001111111111111110111111111111111011;
            32'd15: maze <= 128'b10111111111111111000100000000011111011101111101110001000100000111011101110111111100000100000001111111111111110111111111111111011;
            32'd16: maze <= 128'b10111111111111111010000010000011101110101010111110001010101000111110101011111011100000100000001111111111111110111111111111111011;
            32'd17: maze <= 128'b10111111111111111010000000001011101010111110101110101000101000111011111010111011100000001000001111111111111110111111111111111011;
            32'd18: maze <= 128'b10111111111111111010000000000011101011111111101110100000100000111011111110111011100000000010001111111111111110111111111111111011;
            32'd19: maze <= 128'b10111111111111111000100000100011111011101010111110100010101000111011101010111011100000001000001111111111111110111111111111111011;
            32'd20: maze <= 128'b10111111111111111000001000000011111110101011111110001010100000111011101111111011100000000000001111111111111110111111111111111011;
            32'd21: maze <= 128'b10111111111111111010000000100011101011111010101110101000101010111010101010111011100010100000001111111111111110111111111111111011;
            32'd22: maze <= 128'b10111111111111111010001000001011101010111010101110101000101000111010111010111011100010000010001111111111111110111111111111111011;
            32'd23: maze <= 128'b10111111111111111010000000100011101010111011101110101010101000111011101010101011100000100000101111111111111110111111111111111011;
            32'd24: maze <= 128'b10111111111111111010000000000011101110101111101110001010101000111110111010101111100000001000001111111111111110111111111111111011;
            32'd25: maze <= 128'b10111111111111111010000000001011101011111110101110101000000010111010101111111011100010000000001111111111111110111111111111111011;
            32'd26: maze <= 128'b10111111111111111000001000000011111110101111101110000010101000111011111010101111100000001000001111111111111110111111111111111011;
            32'd27: maze <= 128'b10111111111111111000000000100011111111111011101110001000001000111010101111101011101000000000101111111111111110111111111111111011;
            32'd28: maze <= 128'b10111111111111111010001000000011101010101111101110001000100010111111111110101011100000000010001111111111111110111111111111111011;
            32'd29: maze <= 128'b10111111111111111000001000000011111110111011101110001000101010111011111010101011100000000010001111111111111110111111111111111011;
            32'd30: maze <= 128'b10111111111111111000000000100011111111111010101110100000001010111010111111101011100000000000101111111111111110111111111111111011;
            32'd31: maze <= 128'b10111111111111111010001000100011101010101010101110001010100010111111101011111011100000001000001111111111111110111111111111111011;
            32'd32: maze <= 128'b10111111111111111010001000100011101010101110101110101010000010111010101111111011100010000000001111111111111110111111111111111011;
            32'd33: maze <= 128'b10111111111111111000000000000011111111111111101110000010000010111011101010111011100010001000001111111111111110111111111111111011;
            32'd34: maze <= 128'b10111111111111111000100000100011111010111010101110100010001010111011111011111011100000000000001111111111111110111111111111111011;
            32'd35: maze <= 128'b10111111111111111000000010000011111111101011101110000010101010111011101010101011100010000010001111111111111110111111111111111011;
            32'd36: maze <= 128'b10111111111111111010000010000011101011101011101110101010001010111010101111101011100010000000001111111111111110111111111111111011;
            32'd37: maze <= 128'b10111111111111111010000000100011101011101011101110101000100000111011101111111011100000100000001111111111111110111111111111111011;
            32'd38: maze <= 128'b10111111111111111000000000001011111111111110101110001000001000111011101110111011100000001000001111111111111110111111111111111011;
            32'd39: maze <= 128'b10111111111111111010001000001011101010101010101110001010101000111111101110111011100000000010001111111111111110111111111111111011;
            32'd40: maze <= 128'b10111111111111111010000000100011101011111011101110101000101000111010101110101011100010000000101111111111111110111111111111111011;
            32'd41: maze <= 128'b10111111111111111000000000100011111111111010111110001000101000111010101010111011101000100000001111111111111110111111111111111011;
            32'd42: maze <= 128'b10111111111111111000001000100011111110101010101110001000101010111011111110111011100000000000001111111111111110111111111111111011;
            32'd43: maze <= 128'b10111111111111111010001000001011101010101010101110101000101010111011111110101011100000000010001111111111111110111111111111111011;
            32'd44: maze <= 128'b10111111111111111000000010000011111111101110101110100000100010111010111110111011100000000010001111111111111110111111111111111011;
            32'd45: maze <= 128'b10111111111111111000000010000011111111101011111110100010100000111010101011111011100010000000001111111111111110111111111111111011;
            32'd46: maze <= 128'b10111111111111111000000000100011111111111010101110001000101010111011101010101011100000100000101111111111111110111111111111111011;
            32'd47: maze <= 128'b10111111111111111010000000100011101110111010101110100010001010111010111011101011100010000000101111111111111110111111111111111011;
            32'd48: maze <= 128'b10111111111111111000000000000011111111111111101110000000100010111011111010101011100000100010001111111111111110111111111111111011;
            32'd49: maze <= 128'b10111111111111111010000010001011101010101010101110101010101000111011101010111011100000100010001111111111111110111111111111111011;
            32'd50: maze <= 128'b10111111111111111010000000001011101011111110101110100000101000111011111010111011100000001000001111111111111110111111111111111011;
            32'd51: maze <= 128'b10111111111111111010000000000011101011111111101110100010100000111011101010111111100000100000001111111111111110111111111111111011;
            32'd52: maze <= 128'b10111111111111111010001000000011101010101110101110101000100010111011111110111011100000000010001111111111111110111111111111111011;
            32'd53: maze <= 128'b10111111111111111000000000000011111111111111101110100000000010111010111011111011100000100000001111111111111110111111111111111011;
            32'd54: maze <= 128'b10111111111111111010000000000011101011101111101110100010001010111011111110101011100000000010001111111111111110111111111111111011;
            32'd55: maze <= 128'b10111111111111111000100000100011111011101011101110101000101000111010101110101011100000100000101111111111111110111111111111111011;
            32'd56: maze <= 128'b10111111111111111000100010001011111010101010101110101010001010111010101111101011100000100000001111111111111110111111111111111011;
            32'd57: maze <= 128'b10111111111111111010001000000011101010101011101110101010101010111010101110101011100010000010001111111111111110111111111111111011;
            32'd58: maze <= 128'b10111111111111111010000010000011101110101011101110100010101000111010111011101011100010000000101111111111111110111111111111111011;
            32'd59: maze <= 128'b10111111111111111010000000000011101011111111101110101010000010111010101010111011100010001000001111111111111110111111111111111011;
            32'd60: maze <= 128'b10111111111111111000100000000011111010101111101110101010000010111010111111101011100000000000101111111111111110111111111111111011;
            32'd61: maze <= 128'b10111111111111111000000000000011111111111111101110000000001000111010111111101111101000000000001111111111111110111111111111111011;
            32'd62: maze <= 128'b10111111111111111010000000000011101110111011101110001000101010111110111110101011100000000010001111111111111110111111111111111011;
            32'd63: maze <= 128'b10111111111111111010000000000011101010111111101110101000001000111011111110101111100000000010001111111111111110111111111111111011;
            32'd64: maze <= 128'b10111111111111111000000010000011111111101011101110000010001000111010111111101111101000000000001111111111111110111111111111111011;
            32'd65: maze <= 128'b10111111111111111010000000001011101011101110101110100010001010111011111110101011100000000010001111111111111110111111111111111011;
            32'd66: maze <= 128'b10111111111111111000000010001011111111101010101110100010101010111010101010101011100010000010001111111111111110111111111111111011;
            32'd67: maze <= 128'b10111111111111111000000000001011111111111110101110001000001010111010101110101011101000001000001111111111111110111111111111111011;
            32'd68: maze <= 128'b10111111111111111010000000100011101110111010101110100010001010111010111011111011100010000000001111111111111110111111111111111011;
            32'd69: maze <= 128'b10111111111111111000000000000011111111111111101110100010000010111010101011101011100010000010001111111111111110111111111111111011;
            32'd70: maze <= 128'b10111111111111111010000000000011101011101111101110101000100010111011101110101011100000100010001111111111111110111111111111111011;
            32'd71: maze <= 128'b10111111111111111000000000000011111111111111101110100010000000111010101011111111100010000000001111111111111110111111111111111011;
            32'd72: maze <= 128'b10111111111111111010000000000011101111101111101110100000101000111010111110101111100010000000001111111111111110111111111111111011;
            32'd73: maze <= 128'b10111111111111111000000000001011111111111110101110100010001010111010101010101011100010001000001111111111111110111111111111111011;
            32'd74: maze <= 128'b10111111111111111000001000000011111110101111101110001010001010111010101110101011101000000010001111111111111110111111111111111011;
            32'd75: maze <= 128'b10111111111111111000001000000011111110101110101110000010001010111011111111101011100000000000101111111111111110111111111111111011;
            32'd76: maze <= 128'b10111111111111111000100000000011111010111111101110001000001000111011111111101011100000000000101111111111111110111111111111111011;
            32'd77: maze <= 128'b10111111111111111000100000000011111010111111101110001000100010111011111010101011100000001010001111111111111110111111111111111011;
            32'd78: maze <= 128'b10111111111111111010000000100011101111101010101110000010101010111111101010111011100000001000001111111111111110111111111111111011;
            32'd79: maze <= 128'b10111111111111111000000000000011111111111111101110100000100000111010101110111111100010000000001111111111111110111111111111111011;
            32'd80: maze <= 128'b10111111111111111000100000000011111010111110101110001010001010111011111010111011100000001000001111111111111110111111111111111011;
            32'd81: maze <= 128'b10111111111111111000000010000011111111101010101110000000101010111011111111101011100000000000101111111111111110111111111111111011;
            32'd82: maze <= 128'b10111111111111111010000000000011101111111010101110100000101010111010111011101011100010000000101111111111111110111111111111111011;
            32'd83: maze <= 128'b10111111111111111010000000001011101111111010101110001000101010111110101010101011100000100010001111111111111110111111111111111011;
            32'd84: maze <= 128'b10111111111111111000100000100011111010111010101110001000100010111011111111111011100000000000001111111111111110111111111111111011;
            32'd85: maze <= 128'b10111111111111111010000010001011101011101010101110101010001010111010101111101011100010000000001111111111111110111111111111111011;
            32'd86: maze <= 128'b10111111111111111000000010001011111111101010101110100010101000111010101010111011100010000010001111111111111110111111111111111011;
            32'd87: maze <= 128'b10111111111111111000100000000011111010111111101110001010000000111011101011111111100000100000001111111111111110111111111111111011;
            32'd88: maze <= 128'b10111111111111111010000000000011101011111111101110001000000000111111101111111111100000000000001111111111111110111111111111111011;
            32'd89: maze <= 128'b10111111111111111000100000100011111011101010101110100010100010111011101011111011100000001000001111111111111110111111111111111011;
            32'd90: maze <= 128'b10111111111111111000100000000011111010101111101110001010101000111011111010101111100000001000001111111111111110111111111111111011;
            32'd91: maze <= 128'b10111111111111111010000000100011101011111010101110100000101010111011111010111011100000001000001111111111111110111111111111111011;
            32'd92: maze <= 128'b10111111111111111000000010000011111111101110101110100010001010111010101110101011100010000000101111111111111110111111111111111011;
            32'd93: maze <= 128'b10111111111111111000001000000011111110101111101110001010100010111010101010101011101000001010001111111111111110111111111111111011;
            32'd94: maze <= 128'b10111111111111111000100000000011111011111011101110101000101010111010101010101011100000100010001111111111111110111111111111111011;
            32'd95: maze <= 128'b10111111111111111000000010000011111111101011101110001000101000111010101110101111101000000010001111111111111110111111111111111011;
            32'd96: maze <= 128'b10111111111111111000000010001011111111101010101110100010001000111010101111111011100010000000001111111111111110111111111111111011;
            32'd97: maze <= 128'b10111111111111111000000010001011111111101010101110001000101000111010101110111011101000000010001111111111111110111111111111111011;
            32'd98: maze <= 128'b10111111111111111000000000000011111111111111101110100000001000111010101111101111100010000000001111111111111110111111111111111011;
            32'd99: maze <= 128'b10111111111111111010000000100011101011111011101110101010001000111010101011101011100010000000101111111111111110111111111111111011;
        endcase
    end
    else begin
        maze <= maze;
    end

end
 

endmodule


module CountAndGrade(
    input clk,
    input reset, 
    input end_game,
    output [6:0] out_count_ten,
    output [6:0] out_count,
    output [6:0] out_win_ten,
    output [6:0] out_win,
    output wire refresh_maze
);

wire clk_div;

wire [7:0] count_number;
wire [3:0] count_ten;
wire [3:0] count;

wire [7:0] win_number;
wire [3:0] win_ten;
wire [3:0] win;

wire overtime;

// Instantiate FrequencyDivider module
FrequencyDivider u_FreqDiv (
    .clk(clk),
    .reset(reset),
    .clk_div(clk_div)
);

// Instantiate CounterWithSevenSegment module
CountDownCounter u_count_down (
    .clk(clk_div),
    .reset(reset),
    .refresh_maze(refresh_maze),
    .counter(count_number),
    .overtime(overtime)
);

// Instantiate CalculateGame module
CalculateGame u_cal(
    .clk(clk),
    .reset(reset),
    .end_game(end_game),
    .overtime(overtime),
    .win_counter(win_number),
    .refresh_maze(refresh_maze)
);

// count down counter output to seven seg
NumberToSevenSeg u_num_to_sev0(
    .number(count_number), 
    .out(count), 
    .out_ten(count_ten)
);
SevenSegmentDisplay u_disp0(
    .number(count), 
    .out(out_count)
);
SevenSegmentDisplay u_disp1(
    .number(count_ten), 
    .out(out_count_ten)
);

// win counter output to seven seg
NumberToSevenSeg u_num_to_sev1(
    .number(win_number), 
    .out(win), 
    .out_ten(win_ten)
);
SevenSegmentDisplay u_disp2(
    .number(win), 
    .out(out_win)
);
SevenSegmentDisplay u_disp3(
    .number(win_ten), 
    .out(out_win_ten)
);

endmodule


`define TimeExpire 32'd25000000
module FrequencyDivider (clk,reset,clk_div);
input clk,reset;
output reg clk_div;
reg [31:0] counter_internal;

always @(posedge clk or negedge reset) begin
    if (!reset) begin
        counter_internal <= 32'd0; // Reset the counter
        clk_div <= 1'b0; // Initialize the divided clock
    end else begin
        if (counter_internal == `TimeExpire) begin
            counter_internal <= 32'd0;
            clk_div <= ~clk_div; // Toggle the divided clock
        end else begin
            counter_internal <= counter_internal + 32'd1;
        end
    end
end

endmodule


module NumberToSevenSeg (
    input [7:0] number,
    output reg [6:0] out,
    output reg [6:0] out_ten
);

always @(number)
begin
    out = number % 10;
    out_ten = number / 10;
end

endmodule


module CountDownCounter (
    input wire clk,
    input wire reset,
    input wire refresh_maze,
    output reg [7:0] counter,
    output reg overtime
);

initial begin
    counter = 8'd99;
end

always @(posedge clk or negedge reset or posedge refresh_maze) begin
    if (!reset || refresh_maze) begin
        counter <= 8'd99;
        overtime <= 0;
    end
    else begin
        if (counter == 8'd0) begin
            counter <= 8'd99;
            overtime <= 1;
        end else begin
            counter <= counter - 8'd1;
        end
    end
end


endmodule

module CalculateGame (
    input wire clk,
    input wire reset,
    input wire end_game,
    input wire overtime,
    output reg [7:0] win_counter,
    output reg refresh_maze
);

initial begin
    win_counter = 8'd0;
end

reg [31:0] clk_counter;

always @(posedge clk or negedge reset)begin
    if (!reset) begin
        win_counter <= 8'd0;
        refresh_maze <= 1;
    end else begin
        if (clk_counter == 32'd5000) begin
            clk_counter <= 32'd0;
            if (end_game) begin
                if (!refresh_maze) begin
                    win_counter <= win_counter + 1;
                    refresh_maze <= 1;
                end
            end else if (overtime) begin
                if (!refresh_maze) begin
                    refresh_maze <= 1;
                end
            end else begin
                win_counter <= win_counter;
                refresh_maze <= 0;
            end
        end 
        else begin
            clk_counter <= clk_counter + 1;
        end
    end
end

endmodule

module SevenSegmentDisplay (
    input wire [3:0] number,
    output reg [6:0] out
);

always @(*) begin
    case (number)
        4'b0000: out = 7'b1000000; 
        4'b0001: out = 7'b1111001;
        4'b0010: out = 7'b0100100;
        4'b0011: out = 7'b0110000;
        4'b0100: out = 7'b0011001;
        4'b0101: out = 7'b0010010;
        4'b0110: out = 7'b0000010;
        4'b0111: out = 7'b1111000;
        4'b1000: out = 7'b0000000;
        4'b1001: out = 7'b0010000;
        4'b1010: out = 7'b0001000;
        4'b1011: out = 7'b0000011;
        4'b1100: out = 7'b1000110;
        4'b1101: out = 7'b0100001;
        4'b1110: out = 7'b0000110;
        4'b1111: out = 7'b0001110;
        default: out = 7'b1000000; // 預設輸出為0
    endcase
end

endmodule
 
